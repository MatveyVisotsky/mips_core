library verilog;
use verilog.vl_types.all;
entity insruction_memory_test is
end insruction_memory_test;
